import risc_v_mike_pkg::*;
import UART_MIKE_pkg::*;
//ENDIF
`include "risc_v_mike_header.svh"

module risc_v_mem_ctrl_tb();




endmodule

