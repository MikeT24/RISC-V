module risc_v_mike_top ();

endmodule
